


module XM_datapath 
(
	input wire clk, rst, 

	
);


endmodule
