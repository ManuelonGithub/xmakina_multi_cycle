


module XM_datapath 
(
);


endmodule
