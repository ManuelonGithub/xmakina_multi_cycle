
module bus_interconnect
#(
    parameter WORD = 16,
    parameter SLAVES = 4
 )
(
    input wire[SLAVES-1:0] slaveEn_i, slaveAck_i,
    
);
    

endmodule

